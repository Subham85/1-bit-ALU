* /home/subham109/Downloads/eSim-2.3/library/SubcircuitLibrary/and_gate/and_gate.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 05 Oct 2022 05:18:10 AM PDT

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC1  Net-_SC1-Pad1_ /a /vdd /vdd sky130_fd_pr__pfet_01v8		
SC4  Net-_SC1-Pad1_ /b /vdd /vdd sky130_fd_pr__pfet_01v8		
SC2  Net-_SC1-Pad1_ /a Net-_SC2-Pad3_ Net-_SC2-Pad3_ sky130_fd_pr__nfet_01v8		
SC3  Net-_SC2-Pad3_ /b GND GND sky130_fd_pr__nfet_01v8		
SC5  /y Net-_SC1-Pad1_ /vdd /vdd sky130_fd_pr__pfet_01v8		
SC6  /y Net-_SC1-Pad1_ GND GND sky130_fd_pr__nfet_01v8		
U1  /a /b /vdd /y PORT		

.end
