module fa(input a,b,cin,output reg s,cout);

assign  {cout,s}=a+b+cin;

endmodule
