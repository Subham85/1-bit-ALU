module orgate(input a,b,output c);

or (c,a,b);

endmodule
