* /home/subham109/Downloads/eSim-2.3/library/SubcircuitLibrary/andg/andg.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 05 Oct 2022 06:02:42 AM PDT

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC2  Net-_SC1-Pad1_ /A Net-_SC2-Pad3_ Net-_SC2-Pad3_ sky130_fd_pr__nfet_01v8		
SC1  Net-_SC1-Pad1_ /A /VDD /VDD sky130_fd_pr__pfet_01v8		
SC4  Net-_SC1-Pad1_ /B /VDD /VDD sky130_fd_pr__pfet_01v8		
SC3  Net-_SC2-Pad3_ /B GND GND sky130_fd_pr__nfet_01v8		
U1  /A /B /VDD /Y PORT		
SC5  /Y Net-_SC1-Pad1_ /VDD /VDD sky130_fd_pr__pfet_01v8		
SC6  /Y Net-_SC1-Pad1_ GND GND sky130_fd_pr__nfet_01v8		

.end
